H:\IntelliTank2\intelliTank\schematics\intank.cir
* File created from design "H:\IntelliTank2\intelliTank\schematics\intank.sch" using DesignSpark 17.0.3

U1 +12V GND N0007 L7805CV3 
U2 N0043 unconnected1 N0007 ATMEGA328P-PU 
D1 N0007 N0016 Diode 
CY1 N0016 GND 0.25p Rser=0.1 Lser=0.001 Cpar=5e-011 
XPL1 N0016 N0019 N0020 unconnected2 CONN_SIL_4 
XPL2 N0016 GND N0024 CONN_SIL_3 
Q1 N0028 N0033 GND ZTX450 
Q2 N0029 N0034 GND ZTX450 
Q3 N0030 N0035 GND ZTX450 
R1 N0039 N0030 4k7 
R2 N0040 N0029 4k7 
R3 N0041 N0028 4k7 
XPL3 +12V N0033 N0034 N0035 CONN_SIL_4 
BZ1 GND N0043 ????  
XPL4 N0016 GND N0048 CONN_SIL_3 
XPL5 N0016 GND N0051 CONN_SIL_3 
LDR1 N0016 N0057 ????  
R4 GND N0057 4k7 
LED1 N0065 N0068 LED 3MM GREEN 
LED2 N0060 N0063 LED 3MM RED 
LED3 N0066 N0067 LED 3MM YELLOW 
R5 GND N0063 1K 
R6 GND N0068 1K 
R7 GND N0067 1K 

.tran 0 1m 0 20u
.options Vntol=1u Abstol=1p Reltol=1m
.temp 27



.end
